@00000000
00 00 A0 E3 00 F0 3F E1 00 00 E0 E3 10 0F 03 EE 
01 00 A0 E3 10 0F 02 EE 00 D0 9F E5 42 00 00 EB 
00 40 00 00 1C 30 9F E5 1C 00 9F E5 03 30 60 E0 
06 00 53 E3 0E F0 A0 91 10 30 9F E5 00 00 53 E3 
0E F0 A0 01 03 F0 A0 E1 33 03 00 00 30 03 00 00 
00 00 00 00 24 10 9F E5 24 00 9F E5 01 10 60 E0 
41 11 A0 E1 A1 1F 81 E0 C1 10 B0 E1 0E F0 A0 01 
10 30 9F E5 00 00 53 E3 0E F0 A0 01 03 F0 A0 E1 
30 03 00 00 30 03 00 00 00 00 00 00 10 40 2D E9 
2C 40 9F E5 00 30 D4 E5 00 00 53 E3 06 00 00 1A 
DF FF FF EB 1C 30 9F E5 00 00 53 E3 18 00 9F 15 
00 00 A0 11 01 30 A0 E3 00 30 C4 E5 10 40 BD E8 
0E F0 A0 E1 34 03 00 00 00 00 00 00 30 03 00 00 
40 30 9F E5 00 00 53 E3 10 40 2D E9 38 10 9F 15 
38 00 9F 15 00 00 A0 11 34 00 9F E5 00 30 90 E5 
00 00 53 E3 01 00 00 1A 10 40 BD E8 D4 FF FF EA 
20 30 9F E5 00 00 53 E3 FA FF FF 0A 0F E0 A0 E1 
03 F0 A0 E1 F7 FF FF EA 00 00 00 00 38 03 00 00 
30 03 00 00 2C 03 00 00 00 00 00 00 04 B0 2D E5 
00 B0 8D E2 0C D0 4D E2 1A 3A A0 E3 88 20 A0 E3 
00 20 83 E5 00 30 A0 E3 08 30 0B E5 06 00 00 EA 
1A 3A A0 E3 04 30 83 E2 00 20 A0 E3 00 20 83 E5 
08 30 1B E5 01 30 83 E2 08 30 0B E5 08 30 1B E5 
59 00 53 E3 F5 FF FF DA 1A 3A A0 E3 08 30 83 E2 
C4 20 A0 E3 00 20 83 E5 1A 3A A0 E3 04 30 83 E2 
03 20 A0 E3 00 20 83 E5 00 30 A0 E3 08 30 0B E5 
06 00 00 EA 1A 3A A0 E3 04 30 83 E2 00 20 A0 E3 
00 20 83 E5 08 30 1B E5 01 30 83 E2 08 30 0B E5 
08 30 1B E5 59 00 53 E3 F5 FF FF DA 1A 3A A0 E3 
08 30 83 E2 9E 20 A0 E3 00 20 83 E5 1A 3A A0 E3 
04 30 83 E2 03 20 A0 E3 00 20 83 E5 00 30 A0 E3 
08 30 0B E5 06 00 00 EA 1A 3A A0 E3 04 30 83 E2 
00 20 A0 E3 00 20 83 E5 08 30 1B E5 01 30 83 E2 
08 30 0B E5 08 30 1B E5 59 00 53 E3 F5 FF FF DA 
1A 3A A0 E3 08 30 83 E2 7F 20 A0 E3 00 20 83 E5 
1A 3A A0 E3 04 30 83 E2 03 20 A0 E3 00 20 83 E5 
00 30 A0 E3 08 30 0B E5 06 00 00 EA 1A 3A A0 E3 
04 30 83 E2 00 20 A0 E3 00 20 83 E5 08 30 1B E5 
01 30 83 E2 08 30 0B E5 08 30 1B E5 59 00 53 E3 
F5 FF FF DA 1A 3A A0 E3 08 30 83 E2 70 20 A0 E3 
00 20 83 E5 1A 3A A0 E3 04 30 83 E2 03 20 A0 E3 
00 20 83 E5 00 30 A0 E3 08 30 0B E5 06 00 00 EA 
1A 3A A0 E3 04 30 83 E2 00 20 A0 E3 00 20 83 E5 
08 30 1B E5 01 30 83 E2 08 30 0B E5 08 30 1B E5 
59 00 53 E3 F5 FF FF DA FE FF FF EA 00 00 A0 E3 
00 F0 3F E1 00 00 E0 E3 10 0F 03 EE 01 00 A0 E3 
10 0F 02 EE 00 D0 9F E5 8F FF FF EB 00 40 00 00 
@000002F0
0D C0 A0 E1 F8 DF 2D E9 04 B0 4C E2 28 D0 4B E2 
F0 6F 9D E8 0E F0 A0 E1 
@00000308
0D C0 A0 E1 F8 DF 2D E9 04 B0 4C E2 28 D0 4B E2 
F0 6F 9D E8 0E F0 A0 E1 
@00000320
00 00 00 00 
@00000324
D0 00 00 00 
@00000328
8C 00 00 00 
@0000032C
00 00 00 00 
@00000330
00 00 00 00 
